library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Globals is
    type STATES is (RECEIVING, EDITING, SENDING);
end Globals;

package body Globals is
end Globals;
