library IEEE;
use IEEE.std_logic_1164.all;

package Globals is
    type states is (RECEIVING, EDITING, SENDING);
end Globals;

package body Globals is
end Globals;
